module and_struct(output y,input a,b);
and G1(y,a,b);
endmodule