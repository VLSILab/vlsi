library verilog;
use verilog.vl_types.all;
entity D_ff_tb is
end D_ff_tb;
