module and_gate(y, a, b);
input a;
input b;
output y;
and G1(y, a, b);

endmodule