library verilog;
use verilog.vl_types.all;
entity JK_ff_tb is
end JK_ff_tb;
