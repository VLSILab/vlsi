library verilog;
use verilog.vl_types.all;
entity SR_FF_tb is
end SR_FF_tb;
