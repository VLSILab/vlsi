library verilog;
use verilog.vl_types.all;
entity ParityChecker_tb is
end ParityChecker_tb;
