library verilog;
use verilog.vl_types.all;
entity D_FF_tb is
end D_FF_tb;
