module and_gate(y, a, b);
input a;
input b;
output y;
or G1(y, a, b);

endmodule