library verilog;
use verilog.vl_types.all;
entity tb_async_counter is
end tb_async_counter;
